`timescale 1ns/1ps
module Pipeline_CPU(
    clk_i,
    rst_i
);

//I/O port
input         clk_i;//v
input         rst_i;//v

//myself add
wire [32-1:0] Imm_4 = 4;
wire [32-1:0] instr_o;
wire [32-1:0] zero = 0;
wire [32-1:0] MUX_MemtoReg_out;
wire [1:0] final_mux_select_o;

//Internal Signals
wire [31:0] PC_i; //v
wire [31:0] PC_o; //v
wire [31:0] MUXMemtoReg_o;
wire [31:0] ALUResult;//v
wire [31:0] MUXALUSrc_o;//v
wire [31:0] Decoder_o = {Branch,ALUSrc,RegWrite,ALUOp,MemRead,MemWrite,MemtoReg,Jump};
wire [31:0] RSdata_o;//v
wire [31:0] RTdata_o;//v
wire [31:0] Imm_Gen_o;//v
wire [31:0] ALUSrc1_o;//v
wire [31:0] ALUSrc2_o;//v
wire [31:0]  MUX_control_o;

wire [31:0] PC_Add_Immediate;//v
wire [1:0] ALUOp;//v
wire PC_write;//v
wire ALUSrc;//v
wire RegWrite;//v
wire Branch;//v
wire MUXControl; //v // generated by hazard detection unit
wire Jump;//v
wire [31:0] SL1_o;//v
wire [3:0] ALU_Ctrl_o;//v
wire ALU_zero;//v
wire Branch_zero;
wire MUXPCSrc = ~(Jump|(Branch&ALU_zero));
wire [31:0] DM_o;//v
wire MemtoReg, MemRead, MemWrite;//v
wire [1:0] ForwardA;//v
wire [1:0] ForwardB;//v
wire [31:0] PC_Add4; //v


//Pipeline Register Signals
//IFID
wire [31:0] IFID_PC_o; //v
wire [31:0] IFID_Instr_o;//v
wire IFID_Write; //v
wire IFID_Flush=Branch; //v
wire [31:0]IFID_PC_Add4_o;//v

//IDEXE
wire [31:0] IDEXE_Instr_o;//v
wire [2:0] IDEXE_WB_o; //v
wire [1:0] IDEXE_Mem_o; //v
wire [2:0] IDEXE_Exe_o;//v
wire [31:0] IDEXE_PC_o;
wire [31:0] IDEXE_RSdata_o;//v
wire [31:0] IDEXE_RTdata_o;//v
wire [31:0] IDEXE_ImmGen_o;//v
wire [3:0] IDEXE_Instr_30_14_12_o;//v
wire [4:0] IDEXE_Instr_11_7_o;//v
wire [31:0]IDEXE_PC_add4_o;//v

//EXEMEM
wire [31:0] EXEMEM_Instr_o;//v
wire [2:0] EXEMEM_WB_o;//v
wire [1:0] EXEMEM_Mem_o;//v
wire [31:0] EXEMEM_PCsum_o;
wire EXEMEM_Zero_o;//v
wire [31:0] EXEMEM_ALUResult_o;//v
wire [31:0] EXEMEM_RTdata_o;//v
wire [4:0]  EXEMEM_Instr_11_7_o;//v
wire [31:0] EXEMEM_PC_Add4_o; //v

//MEMWB
wire [2:0] MEMWB_WB_o;//v
wire [31:0] MEMWB_DM_o;//v
wire [31:0] MEMWB_ALUresult_o;//v
wire [4:0]  MEMWB_Instr_11_7_o;//v
wire [31:0] MEMWB_PC_Add4_o;//v


// IF
MUX_2to1 MUX_PCSrc(
    PC_Add_Immediate,//data1
    PC_Add4,
    MUXPCSrc,//select
    PC_i
);

ProgramCounter PC(
    clk_i,
    rst_i,
    PC_write,
    PC_i,
    PC_o
);

Adder PC_plus_4_Adder(
    PC_o,
    Imm_4,
    PC_Add4
);

Instr_Memory IM(
    PC_o,
    instr_o
);

IFID_register IFtoID(  
    clk_i,
    rst_i,
    IFID_Write,
    IFID_Flush,
    PC_o,
    instr_o,
    PC_Add4,
    IFID_PC_o,
    IFID_Instr_o,
    IFID_PC_Add4_o
);

// ID
Hazard_detection Hazard_detection_obj(
    IFID_Instr_o[19:15],//ifid_regrs
    IFID_Instr_o[24:20],//ifid_regrt
    IDEXE_Instr_11_7_o,//idexe_regrd
    IDEXE_Mem_o[1],//idexe_memread
    PC_write,//pc_write
    IFID_Write,//ifid_write
    MUXControl//control_output_select
);

MUX_2to1 MUX_control( //?
    Decoder_o,//data1
    zero,//data2
    MUXControl,//select
    MUX_control_o//output
);

Decoder Decoder(
    IFID_Instr_o,//instri
    Branch,//branch
    ALUSrc,//alusrc
    RegWrite,//regwrite
    ALUOp,//aluop
    MemRead,//memread
    MemWrite,//memwrite
    MemtoReg,//memtoreg
    Jump//jump
);

Reg_File RF(
    clk_i,//clk
    rst_i,//rst
    IFID_Instr_o[19:15],//rsaddri
    IFID_Instr_o[24:20],//rtaddri
    MEMWB_Instr_11_7_o,//rdaddri
    MUX_MemtoReg_out,//rdatati
    MEMWB_WB_o[1],//regwritei
    RSdata_o,//rsdatao
    RTdata_o//rtdatao
);

Imm_Gen ImmGen(
    IFID_Instr_o,//instri
    Imm_Gen_o//imm_gen_o
);

Shift_Left_1 SL1(
    Imm_Gen_o,//datai
    SL1_o//datao
);

Adder Branch_Adder(
    SL1_o,//src1
    IFID_PC_o,//src2
    PC_Add_Immediate//sum
);

IDEXE_register IDtoEXE(
    clk_i,//clk
    rst_i,//rst
    IFID_Instr_o,//instri
    {Jump,RegWrite,MemtoReg},//wbi
    {MemRead,MemWrite},//memi
    {ALUOp,ALUSrc},//exei
    RSdata_o,//data1i
    RTdata_o,//data2i
    Imm_Gen_o,//immgeni
    {IFID_Instr_o[30],IFID_Instr_o[14:12]},//aluctrl_instr
    IFID_Instr_o[11:7],//wbregi
    IFID_PC_Add4_o,//pc_add4_i
    IDEXE_Instr_o,//instro
    IDEXE_WB_o,//wbo
    IDEXE_Mem_o,//memo
    IDEXE_Exe_o,//exeo
    IDEXE_RSdata_o,//data1o
    IDEXE_RTdata_o,//data2o
    IDEXE_ImmGen_o,//immgeno
    IDEXE_Instr_30_14_12_o,//aluctrlinput
    IDEXE_Instr_11_7_o,//wbrego
    IDEXE_PC_add4_o//pcadd4o
);

// EXE
MUX_2to1 MUX_ALUSrc(
    ALUSrc2_o,//data1
    IDEXE_ImmGen_o,//data2
    IDEXE_Exe_o[0],//select
    MUXALUSrc_o//output
);

ForwardingUnit FWUnit(
    IDEXE_Instr_o[19:15],//id_exe_rs1
    IDEXE_Instr_o[24:20],//id_exe_rs2
    EXEMEM_Instr_11_7_o,//exemem_rd
    MEMWB_Instr_11_7_o,//memwb_rd
    EXEMEM_WB_o[1],//exemem_regwrite
    MEMWB_WB_o[1],//memwb_regwrite
    ForwardA,//forwarda
    ForwardB//forwardb
);

MUX_3to1 MUX_ALU_src1(
    IDEXE_RSdata_o,//data0_i,
    MUX_MemtoReg_out,//data1_i,
    EXEMEM_ALUResult_o,//data2_i,
    ForwardA,//select_i,
    ALUSrc1_o//data_o
);

MUX_3to1 MUX_ALU_src2(
    IDEXE_RTdata_o,//data0_i,
    MUX_MemtoReg_out,//data1_i,
    EXEMEM_ALUResult_o,//data2_i,
    ForwardB,//select_i,
    ALUSrc2_o//data_o
);

ALU_Ctrl ALU_Ctrl(
    IDEXE_Instr_30_14_12_o,//instr,
    IDEXE_Exe_o[2:1],//ALUOp,
    ALU_Ctrl_o//ALU_Ctrl_o
);

alu alu(
    rst_i,//rst_n,      
    ALUSrc1_o,//src1,       
    MUXALUSrc_o,//src2,       
    ALU_Ctrl_o,//ALU_control,
    ALUResult,//result,     
    ALU_zero//zero
);

EXEMEM_register EXEtoMEM(
    clk_i,//clk_i,
    rst_i,//rst_i,
    IDEXE_Instr_o,// instr_i,
    IDEXE_WB_o,//WB_i,
    IDEXE_Mem_o,//Mem_i,
    ALU_zero,//zero_i,
    ALUResult,// alu_ans_i,
    IDEXE_RTdata_o,// rtdata_i,
    IDEXE_Instr_11_7_o,//WBreg_i,
    IDEXE_PC_add4_o,// pc_add4_i,

    EXEMEM_Instr_o,// instr_o,
    EXEMEM_WB_o,//WB_o,
    EXEMEM_Mem_o,//Mem_o,
    EXEMEM_Zero_o,//zero_o,
    EXEMEM_ALUResult_o,// alu_ans_o,
    EXEMEM_RTdata_o,// rtdata_o,
    EXEMEM_Instr_11_7_o,//WBreg_o,
    EXEMEM_PC_Add4_o// pc_add4_o
);

// MEM
Data_Memory Data_Memory(
    clk_i,//clk_i,
    EXEMEM_ALUResult_o,//addr_i,
    EXEMEM_RTdata_o,//data_i,
    EXEMEM_Mem_o[1],//MemRead_i,
    EXEMEM_Mem_o[0],//MemWrite_i,
    DM_o//data_o
);

MEMWB_register MEMtoWB(
    clk_i,//clk_i,
    rst_i,//rst_i,
    EXEMEM_WB_o,//WB_i,
    DM_o,// DM_i,
    EXEMEM_ALUResult_o,// alu_ans_i,
    EXEMEM_Instr_11_7_o,//WBreg_i,
    EXEMEM_PC_Add4_o,// pc_add4_i,
    MEMWB_WB_o,//WB_o,
    MEMWB_DM_o,// DM_o,
    MEMWB_ALUresult_o,// alu_ans_o,
    MEMWB_Instr_11_7_o,//WBreg_o,
    MEMWB_PC_Add4_o// pc_add4_o
);

Generate_final_mux_select final_mux_select(
    MEMWB_WB_o[2],
    MEMWB_WB_o[1],
    MEMWB_WB_o[0],
    final_mux_select_o
);
// WB
MUX_3to1 MUX_MemtoReg(
    MEMWB_DM_o,//data0_i,
    MEMWB_ALUresult_o,//data1_i,
    MEMWB_PC_Add4_o,//data2_i,
    final_mux_select_o,//select_i,
    MUX_MemtoReg_out//data_o
);

endmodule
